
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.gfx_util_pkg.all;

package bb_rom_pkg is

	constant MEMORY_CONTENTS : bb_rom_t(0 to 16383) := (
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"7", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"0", x"0", x"0", x"9", x"9", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"b", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"3", x"0", x"0", x"0", x"0", x"9", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"8", x"4", x"4", x"7", x"d", x"f", x"f", x"f", x"f", x"8", x"0", x"0", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"b", x"b", x"0", x"0", x"7", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"6", x"3", x"6", x"a", x"f", x"f", x"f", x"f", x"1", x"1", x"1", x"1", x"e", x"e", x"e", x"e",
	x"f", x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"8", x"0", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"9", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"0", x"0", x"1", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"7", x"0", x"0", x"0", x"0", x"7", x"d", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"8", x"f", x"f", x"f", x"1", x"1", x"1", x"1", x"e", x"e", x"e", x"e",
	x"f", x"f", x"b", x"0", x"0", x"7", x"7", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"a", x"c", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"d", x"9", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"d", x"1", x"0", x"6", x"c", x"d", x"c", x"f", x"f", x"f", x"f", x"f", x"8", x"8", x"9", x"d", x"8", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"8", x"0", x"2", x"e", x"9", x"0", x"0", x"d", x"f", x"f", x"2", x"2", x"2", x"2", x"d", x"d", x"d", x"d",
	x"f", x"f", x"b", x"0", x"0", x"b", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"7", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"9", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"5", x"9", x"f", x"f", x"f", x"f", x"f", x"f", x"b", x"0", x"0", x"7", x"6", x"6", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"8", x"f", x"f", x"f", x"f", x"f", x"b", x"0", x"0", x"7", x"7", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"7", x"0", x"2", x"d", x"9", x"0", x"0", x"b", x"f", x"f", x"2", x"2", x"2", x"2", x"d", x"d", x"d", x"d",
	x"f", x"f", x"b", x"0", x"0", x"d", x"d", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"6", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"9", x"9", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"6", x"f", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"8", x"0", x"0", x"8", x"f", x"f", x"f", x"f", x"f", x"f", x"7", x"0", x"0", x"0", x"0", x"7", x"d", x"f", x"f", x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"3", x"3", x"3", x"3", x"c", x"c", x"c", x"c",
	x"f", x"f", x"b", x"0", x"0", x"b", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"6", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"b", x"3", x"0", x"0", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"d", x"6", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"b", x"b", x"0", x"0", x"8", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"8", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"b", x"b", x"0", x"0", x"9", x"f", x"f", x"f", x"f", x"f", x"a", x"5", x"6", x"7", x"0", x"0", x"c", x"f", x"f", x"3", x"3", x"3", x"3", x"c", x"c", x"c", x"c",
	x"f", x"f", x"b", x"0", x"0", x"7", x"7", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"6", x"0", x"0", x"8", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"9", x"c", x"c", x"3", x"0", x"0", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"d", x"8", x"c", x"c", x"5", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"b", x"0", x"0", x"9", x"f", x"f", x"f", x"f", x"f", x"f", x"8", x"0", x"0", x"8", x"f", x"f", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"b", x"b", x"0", x"0", x"8", x"f", x"f", x"f", x"f", x"f", x"c", x"d", x"c", x"5", x"0", x"0", x"f", x"f", x"f", x"4", x"4", x"4", x"4", x"b", x"b", x"b", x"b",
	x"f", x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"8", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"f", x"d", x"d", x"d", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"8", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"8", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"8", x"d", x"f", x"f", x"f", x"f", x"f", x"f", x"8", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"8", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"4", x"4", x"4", x"4", x"b", x"b", x"b", x"b",
	x"f", x"f", x"f", x"f", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"b", x"8", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"b", x"8", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"b", x"8", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"6", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"b", x"8", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"b", x"8", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"5", x"5", x"5", x"5", x"a", x"a", x"a", x"a",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"5", x"5", x"5", x"5", x"a", x"a", x"a", x"a",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"6", x"6", x"6", x"6", x"9", x"9", x"9", x"9",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"6", x"6", x"6", x"6", x"9", x"9", x"9", x"9",
	x"f", x"f", x"f", x"b", x"0", x"0", x"4", x"f", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"1", x"5", x"8", x"d", x"f", x"f", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"d", x"f", x"f", x"7", x"7", x"7", x"7", x"8", x"8", x"8", x"8",
	x"f", x"f", x"f", x"4", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"3", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"c", x"2", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"d", x"f", x"7", x"7", x"7", x"7", x"8", x"8", x"8", x"8",
	x"f", x"f", x"c", x"0", x"0", x"1", x"0", x"6", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"7", x"d", x"d", x"3", x"0", x"0", x"f", x"f", x"f", x"f", x"4", x"0", x"0", x"7", x"a", x"8", x"0", x"0", x"0", x"f", x"f", x"d", x"0", x"0", x"5", x"b", x"b", x"6", x"0", x"0", x"c", x"f", x"f", x"d", x"0", x"0", x"6", x"c", x"c", x"c", x"c", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"6", x"c", x"c", x"c", x"c", x"f", x"f", x"f", x"f", x"f", x"4", x"0", x"0", x"7", x"a", x"8", x"8", x"0", x"0", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"d", x"f", x"8", x"8", x"8", x"8", x"7", x"7", x"7", x"7",
	x"f", x"f", x"6", x"0", x"4", x"a", x"0", x"0", x"d", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"b", x"0", x"0", x"7", x"f", x"f", x"f", x"d", x"d", x"d", x"f", x"f", x"d", x"0", x"0", x"7", x"f", x"f", x"e", x"4", x"0", x"0", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"c", x"f", x"f", x"d", x"0", x"0", x"6", x"c", x"c", x"c", x"e", x"f", x"f", x"f", x"f", x"b", x"0", x"0", x"7", x"f", x"f", x"f", x"d", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"d", x"f", x"8", x"8", x"8", x"8", x"7", x"7", x"7", x"7",
	x"f", x"d", x"0", x"0", x"a", x"e", x"1", x"0", x"8", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"7", x"f", x"f", x"f", x"a", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"7", x"f", x"f", x"f", x"7", x"0", x"0", x"c", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"c", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"c", x"f", x"f", x"a", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"d", x"f", x"9", x"9", x"9", x"9", x"6", x"6", x"6", x"6",
	x"f", x"8", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"d", x"0", x"0", x"7", x"e", x"e", x"9", x"0", x"0", x"b", x"f", x"f", x"b", x"0", x"0", x"7", x"f", x"f", x"f", x"d", x"d", x"d", x"f", x"f", x"d", x"0", x"0", x"7", x"f", x"f", x"e", x"4", x"0", x"0", x"f", x"f", x"d", x"0", x"0", x"7", x"d", x"d", x"d", x"f", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"c", x"f", x"f", x"b", x"0", x"0", x"7", x"f", x"f", x"f", x"d", x"0", x"0", x"f", x"f", x"c", x"0", x"0", x"4", x"c", x"c", x"c", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"d", x"f", x"9", x"9", x"9", x"9", x"6", x"6", x"6", x"6",
	x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"9", x"f", x"f", x"d", x"0", x"0", x"7", x"e", x"d", x"8", x"0", x"0", x"9", x"f", x"f", x"f", x"4", x"0", x"0", x"7", x"a", x"8", x"0", x"0", x"0", x"f", x"f", x"d", x"0", x"0", x"5", x"c", x"b", x"6", x"0", x"0", x"6", x"f", x"f", x"d", x"0", x"0", x"6", x"c", x"c", x"c", x"c", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"4", x"0", x"0", x"7", x"a", x"8", x"0", x"0", x"0", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"b", x"b", x"b", x"b", x"0", x"0", x"d", x"f", x"a", x"a", x"a", x"a", x"5", x"5", x"5", x"5",
	x"a", x"0", x"0", x"b", x"d", x"d", x"d", x"4", x"0", x"2", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"9", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"3", x"e", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"d", x"0", x"0", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"2", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"d", x"f", x"a", x"a", x"a", x"a", x"5", x"5", x"5", x"5",
	x"a", x"0", x"2", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"b", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"4", x"7", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"0", x"0", x"9", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"d", x"0", x"0", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"0", x"0", x"f", x"0", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"b", x"b", x"b", x"b", x"4", x"4", x"4", x"4",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"b", x"b", x"b", x"b", x"4", x"4", x"4", x"4",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"c", x"c", x"c", x"3", x"3", x"3", x"3",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"c", x"c", x"c", x"3", x"3", x"3", x"3",
	x"c", x"0", x"0", x"b", x"f", x"d", x"d", x"0", x"0", x"0", x"b", x"f", x"f", x"c", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"9", x"f", x"f", x"f", x"f", x"f", x"d", x"8", x"0", x"0", x"0", x"8", x"c", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"9", x"f", x"f", x"f", x"f", x"d", x"0", x"1", x"1", x"1", x"1", x"1", x"1", x"a", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"d", x"d", x"d", x"d", x"2", x"2", x"2", x"2",
	x"c", x"0", x"0", x"b", x"f", x"d", x"0", x"0", x"0", x"b", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"6", x"f", x"f", x"f", x"6", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"0", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"f", x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"9", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"1", x"1", x"0", x"1", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"d", x"d", x"d", x"d", x"2", x"2", x"2", x"2",
	x"c", x"0", x"0", x"a", x"d", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"b", x"f", x"b", x"0", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"0", x"b", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"0", x"0", x"3", x"b", x"b", x"b", x"5", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"a", x"a", x"d", x"d", x"0", x"0", x"0", x"c", x"f", x"f", x"2", x"0", x"4", x"b", x"c", x"c", x"5", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"a", x"a", x"d", x"d", x"0", x"0", x"0", x"c", x"f", x"a", x"0", x"0", x"b", x"c", x"c", x"c", x"c", x"c", x"c", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"1", x"1", x"1", x"1",
	x"c", x"0", x"0", x"2", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"4", x"f", x"4", x"0", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"0", x"0", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"b", x"0", x"0", x"b", x"f", x"c", x"0", x"0", x"b", x"b", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"d", x"0", x"0", x"9", x"f", x"c", x"0", x"0", x"b", x"b", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"9", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"1", x"1", x"1", x"1",
	x"c", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"9", x"0", x"0", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"c", x"c", x"0", x"0", x"c", x"f", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"b", x"0", x"0", x"b", x"f", x"c", x"0", x"0", x"a", x"a", x"d", x"d", x"0", x"0", x"0", x"c", x"f", x"9", x"0", x"0", x"d", x"f", x"f", x"f", x"e", x"0", x"0", x"7", x"f", x"c", x"0", x"0", x"a", x"a", x"d", x"d", x"0", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0",
	x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"8", x"0", x"0", x"0", x"8", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"8", x"0", x"0", x"0", x"c", x"0", x"0", x"c", x"f", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"b", x"0", x"0", x"b", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"b", x"0", x"0", x"b", x"f", x"f", x"f", x"d", x"0", x"0", x"9", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"e", x"9", x"c", x"c", x"c", x"c", x"d", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0",
	x"c", x"0", x"0", x"b", x"b", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"a", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"0", x"0", x"0", x"c", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"c", x"c", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"0", x"0", x"4", x"b", x"b", x"b", x"5", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"1", x"0", x"3", x"b", x"b", x"b", x"5", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"a", x"c", x"c", x"c", x"c", x"c", x"b", x"0", x"0", x"9", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"0", x"0", x"b", x"f", x"b", x"0", x"0", x"0", x"0", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"d", x"c", x"0", x"c", x"d", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"d", x"c", x"c", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"9", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"9", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"a", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"0", x"0", x"b", x"f", x"e", x"b", x"b", x"0", x"0", x"b", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"c", x"0", x"0", x"d", x"f", x"d", x"f", x"d", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"d", x"f", x"d", x"c", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"0", x"0", x"0", x"c", x"f", x"d", x"9", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"c", x"0", x"0", x"0", x"6", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"0", x"0", x"7", x"f", x"f", x"2", x"0", x"3", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"c", x"0", x"0", x"e", x"f", x"f", x"f", x"e", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"0", x"0", x"7", x"f", x"f", x"9", x"0", x"0", x"c", x"f", x"f", x"8", x"0", x"2", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"b", x"0", x"0", x"c", x"f", x"f", x"0", x"0", x"0", x"c", x"c", x"c", x"0", x"0", x"0", x"f", x"f", x"f", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"0", x"0", x"0", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"c", x"c", x"c", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"0", x"0", x"7", x"f", x"f", x"d", x"0", x"0", x"7", x"f", x"f", x"1", x"0", x"9", x"f", x"f", x"c", x"0", x"0", x"b", x"f", x"0", x"f", x"b", x"0", x"0", x"c", x"f", x"f", x"f", x"0", x"0", x"0", x"c", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"c", x"c", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"d", x"d", x"c", x"c", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"0", x"0", x"7", x"f", x"f", x"f", x"6", x"0", x"0", x"e", x"b", x"0", x"0", x"d", x"f", x"f", x"c", x"0", x"0", x"b", x"0", x"0", x"0", x"b", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"0", x"0", x"7", x"f", x"f", x"f", x"b", x"0", x"0", x"a", x"5", x"0", x"6", x"f", x"f", x"f", x"c", x"0", x"0", x"b", x"0", x"0", x"0", x"b", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"a", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"c", x"c", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"0", x"0", x"a", x"f", x"f", x"f", x"f", x"0", x"0", x"8", x"f", x"f", x"f", x"f", x"2", x"0", x"2", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"0", x"0", x"0", x"b", x"b", x"b", x"0", x"0", x"0", x"b", x"f", x"f", x"f", x"f", x"9", x"0", x"0", x"0", x"2", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"c", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"c", x"d", x"d", x"d", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"9", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"f", x"f", x"f", x"f", x"f", x"d", x"0", x"0", x"0", x"9", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"f", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"c", x"f", x"c", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"c", x"c", x"c", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"b", x"0", x"0", x"0", x"0", x"0", x"9", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"5", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"f", x"0", x"0", x"c", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"b", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"c", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"c", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"3", x"3", x"0", x"0", x"0", x"0", x"0", x"0", x"3", x"3", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"5", x"7", x"7", x"7", x"7", x"6", x"6", x"7", x"7", x"6", x"2", x"6", x"b", x"b", x"8", x"9", x"8", x"8", x"9", x"8", x"b", x"b", x"6", x"3", x"3", x"0", x"7", x"7", x"0", x"0", x"7", x"7", x"0", x"3", x"3", x"0", x"c", x"c", x"c", x"c", x"c", x"c", x"c", x"c", x"c", x"c", x"0", x"3", x"5", x"5", x"4", x"5", x"5", x"5", x"5", x"4", x"5", x"5", x"3", x"0", x"c", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"c", x"0", x"5", x"5", x"5", x"7", x"5", x"5", x"5", x"5", x"7", x"5", x"5", x"5", x"7", x"e", x"d", x"d", x"d", x"0", x"0", x"d", x"d", x"d", x"e", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"6", x"9", x"a", x"a", x"a", x"9", x"a", x"a", x"8", x"6", x"2", x"6", x"a", x"9", x"3", x"5", x"8", x"8", x"5", x"3", x"9", x"a", x"6", x"3", x"0", x"7", x"7", x"0", x"b", x"b", x"0", x"7", x"7", x"0", x"3", x"0", x"c", x"b", x"b", x"b", x"b", x"b", x"b", x"b", x"b", x"c", x"0", x"3", x"5", x"5", x"6", x"5", x"5", x"5", x"5", x"6", x"5", x"5", x"3", x"0", x"5", x"c", x"c", x"3", x"3", x"3", x"3", x"c", x"c", x"5", x"0", x"5", x"7", x"5", x"7", x"5", x"0", x"0", x"5", x"7", x"5", x"7", x"5", x"7", x"d", x"c", x"f", x"3", x"1", x"1", x"3", x"f", x"c", x"d", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"7", x"9", x"9", x"a", x"b", x"b", x"b", x"a", x"8", x"6", x"2", x"6", x"9", x"6", x"1", x"3", x"7", x"7", x"3", x"1", x"6", x"9", x"6", x"0", x"7", x"7", x"0", x"b", x"b", x"b", x"b", x"0", x"7", x"7", x"0", x"0", x"c", x"b", x"0", x"0", x"0", x"0", x"0", x"0", x"b", x"c", x"0", x"3", x"5", x"6", x"5", x"6", x"3", x"3", x"6", x"5", x"6", x"5", x"3", x"0", x"5", x"c", x"c", x"3", x"3", x"3", x"3", x"c", x"c", x"5", x"0", x"5", x"7", x"5", x"5", x"5", x"0", x"0", x"5", x"5", x"5", x"7", x"5", x"7", x"b", x"e", x"2", x"1", x"5", x"5", x"1", x"2", x"e", x"b", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"6", x"9", x"b", x"b", x"b", x"b", x"b", x"b", x"a", x"7", x"2", x"6", x"a", x"7", x"4", x"6", x"8", x"8", x"6", x"4", x"7", x"a", x"6", x"0", x"7", x"0", x"b", x"b", x"0", x"0", x"b", x"b", x"0", x"7", x"0", x"0", x"c", x"b", x"0", x"3", x"3", x"3", x"3", x"0", x"b", x"c", x"0", x"3", x"5", x"5", x"5", x"3", x"c", x"c", x"3", x"5", x"5", x"5", x"3", x"0", x"5", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"5", x"0", x"5", x"7", x"7", x"5", x"0", x"0", x"0", x"0", x"5", x"7", x"7", x"5", x"7", x"f", x"3", x"0", x"3", x"5", x"5", x"3", x"0", x"3", x"f", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"5", x"8", x"a", x"b", x"a", x"9", x"a", x"b", x"a", x"7", x"2", x"6", x"a", x"a", x"9", x"9", x"8", x"8", x"9", x"9", x"a", x"a", x"6", x"0", x"0", x"b", x"b", x"0", x"b", x"b", x"0", x"b", x"b", x"0", x"0", x"0", x"c", x"b", x"0", x"3", x"3", x"3", x"3", x"0", x"b", x"c", x"0", x"3", x"5", x"5", x"3", x"c", x"c", x"c", x"c", x"3", x"5", x"5", x"3", x"0", x"5", x"3", x"3", x"3", x"c", x"c", x"3", x"3", x"3", x"5", x"0", x"5", x"0", x"7", x"5", x"0", x"5", x"5", x"0", x"5", x"7", x"0", x"5", x"7", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"6", x"9", x"b", x"b", x"b", x"a", x"a", x"a", x"8", x"6", x"2", x"6", x"a", x"a", x"9", x"9", x"8", x"8", x"9", x"9", x"a", x"a", x"6", x"0", x"0", x"b", x"b", x"0", x"b", x"b", x"0", x"b", x"b", x"0", x"0", x"0", x"c", x"b", x"0", x"3", x"3", x"3", x"3", x"0", x"b", x"c", x"0", x"3", x"5", x"5", x"3", x"c", x"c", x"c", x"c", x"3", x"5", x"5", x"3", x"0", x"5", x"3", x"3", x"3", x"c", x"c", x"3", x"3", x"3", x"5", x"0", x"0", x"5", x"7", x"0", x"5", x"0", x"0", x"5", x"0", x"7", x"5", x"0", x"7", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"7", x"9", x"a", x"a", x"b", x"a", x"a", x"a", x"9", x"6", x"2", x"6", x"a", x"7", x"4", x"6", x"8", x"8", x"6", x"4", x"7", x"a", x"6", x"0", x"7", x"0", x"b", x"b", x"0", x"0", x"b", x"b", x"0", x"7", x"0", x"0", x"c", x"b", x"0", x"3", x"3", x"3", x"3", x"0", x"b", x"c", x"0", x"3", x"5", x"5", x"5", x"3", x"c", x"c", x"3", x"5", x"5", x"5", x"3", x"0", x"5", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"5", x"0", x"0", x"7", x"7", x"0", x"5", x"5", x"5", x"5", x"0", x"7", x"7", x"0", x"7", x"f", x"3", x"0", x"3", x"5", x"5", x"3", x"0", x"3", x"f", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"7", x"9", x"a", x"a", x"a", x"a", x"a", x"b", x"a", x"7", x"2", x"6", x"9", x"6", x"1", x"3", x"7", x"7", x"3", x"1", x"6", x"9", x"6", x"0", x"7", x"7", x"0", x"b", x"b", x"b", x"b", x"0", x"7", x"7", x"0", x"0", x"c", x"b", x"0", x"0", x"0", x"0", x"0", x"0", x"b", x"c", x"0", x"3", x"5", x"6", x"5", x"6", x"3", x"3", x"6", x"5", x"6", x"5", x"3", x"0", x"5", x"c", x"c", x"3", x"3", x"3", x"3", x"c", x"c", x"5", x"0", x"0", x"7", x"0", x"0", x"0", x"5", x"5", x"0", x"0", x"0", x"7", x"0", x"7", x"b", x"e", x"2", x"1", x"5", x"5", x"1", x"2", x"e", x"b", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"7", x"a", x"b", x"a", x"a", x"b", x"b", x"a", x"9", x"7", x"2", x"6", x"a", x"9", x"3", x"5", x"8", x"8", x"5", x"3", x"9", x"a", x"6", x"3", x"0", x"7", x"7", x"0", x"b", x"b", x"0", x"7", x"7", x"0", x"3", x"0", x"c", x"b", x"b", x"b", x"b", x"b", x"b", x"b", x"b", x"c", x"0", x"3", x"5", x"5", x"6", x"5", x"5", x"5", x"5", x"6", x"5", x"5", x"3", x"0", x"5", x"c", x"c", x"3", x"3", x"3", x"3", x"c", x"c", x"5", x"0", x"0", x"7", x"0", x"7", x"0", x"5", x"5", x"0", x"7", x"0", x"7", x"0", x"7", x"d", x"c", x"f", x"3", x"1", x"1", x"3", x"f", x"c", x"d", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"6", x"9", x"b", x"a", x"9", x"a", x"b", x"a", x"8", x"6", x"2", x"6", x"b", x"b", x"8", x"9", x"8", x"8", x"9", x"8", x"b", x"b", x"6", x"3", x"3", x"0", x"7", x"7", x"0", x"0", x"7", x"7", x"0", x"3", x"3", x"0", x"c", x"c", x"c", x"c", x"c", x"c", x"c", x"c", x"c", x"c", x"0", x"3", x"5", x"5", x"4", x"5", x"5", x"5", x"5", x"4", x"5", x"5", x"3", x"0", x"c", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"c", x"0", x"0", x"0", x"0", x"7", x"0", x"0", x"0", x"0", x"7", x"0", x"0", x"0", x"7", x"e", x"d", x"d", x"d", x"0", x"0", x"d", x"d", x"d", x"e", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"2", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"3", x"3", x"0", x"0", x"0", x"0", x"0", x"0", x"3", x"3", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"7", x"7", x"7", x"0", x"7", x"7", x"7", x"6", x"6", x"0", x"7", x"a", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"6", x"6", x"7", x"0", x"7", x"6", x"6", x"6", x"6", x"0", x"7", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"e", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"c", x"a", x"a", x"c", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"7", x"7", x"6", x"6", x"6", x"0", x"7", x"7", x"6", x"6", x"6", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"9", x"4", x"5", x"9", x"d", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"7", x"7", x"7", x"6", x"6", x"0", x"7", x"7", x"7", x"6", x"6", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"e", x"e", x"e", x"d", x"d", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"e", x"c", x"6", x"0", x"2", x"7", x"c", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"7", x"6", x"7", x"6", x"6", x"0", x"7", x"6", x"7", x"6", x"6", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"d", x"c", x"b", x"a", x"9", x"8", x"9", x"b", x"e", x"f", x"f", x"f", x"f", x"e", x"e", x"a", x"4", x"1", x"2", x"6", x"b", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"b", x"9", x"7", x"5", x"3", x"2", x"2", x"5", x"a", x"e", x"e", x"f", x"f", x"f", x"e", x"d", x"9", x"5", x"5", x"4", x"3", x"9", x"d", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"6", x"0", x"7", x"7", x"6", x"6", x"6", x"0", x"7", x"7", x"6", x"6", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"e", x"e", x"e", x"e", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"a", x"6", x"3", x"3", x"3", x"5", x"5", x"2", x"4", x"a", x"e", x"e", x"f", x"f", x"f", x"e", x"c", x"8", x"7", x"8", x"6", x"1", x"7", x"c", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"6", x"0", x"7", x"7", x"7", x"6", x"6", x"0", x"7", x"7", x"7", x"6", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"e", x"e", x"d", x"d", x"c", x"b", x"b", x"a", x"b", x"c", x"d", x"e", x"e", x"f", x"f", x"f", x"f", x"e", x"d", x"a", x"5", x"3", x"5", x"8", x"a", x"b", x"a", x"5", x"4", x"a", x"e", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"8", x"a", x"8", x"2", x"6", x"b", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"6", x"0", x"7", x"6", x"7", x"6", x"6", x"0", x"7", x"6", x"7", x"6", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"c", x"b", x"a", x"9", x"8", x"6", x"5", x"4", x"4", x"5", x"7", x"a", x"d", x"e", x"f", x"f", x"f", x"e", x"e", x"b", x"6", x"2", x"5", x"9", x"c", x"e", x"e", x"c", x"7", x"5", x"a", x"e", x"f", x"f", x"f", x"e", x"e", x"a", x"6", x"a", x"c", x"9", x"4", x"4", x"a", x"d", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"e", x"c", x"8", x"5", x"4", x"3", x"2", x"3", x"4", x"4", x"2", x"1", x"1", x"4", x"9", x"d", x"e", x"f", x"f", x"e", x"c", x"8", x"2", x"4", x"9", x"d", x"e", x"f", x"f", x"d", x"a", x"a", x"c", x"e", x"f", x"f", x"f", x"e", x"d", x"8", x"6", x"b", x"d", x"b", x"5", x"2", x"8", x"c", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"7", x"7", x"7", x"0", x"7", x"7", x"7", x"6", x"6", x"0", x"7", x"7", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"e", x"e", x"e", x"d", x"d", x"d", x"d", x"d", x"e", x"e", x"f", x"f", x"e", x"b", x"5", x"1", x"0", x"1", x"5", x"8", x"a", x"9", x"8", x"5", x"2", x"1", x"6", x"b", x"e", x"f", x"f", x"e", x"a", x"5", x"1", x"7", x"c", x"e", x"f", x"f", x"f", x"e", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"e", x"c", x"7", x"7", x"c", x"e", x"c", x"6", x"0", x"6", x"b", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"d", x"d", x"c", x"b", x"a", x"9", x"8", x"7", x"8", x"9", x"b", x"d", x"e", x"f", x"e", x"c", x"9", x"6", x"2", x"2", x"8", x"c", x"d", x"d", x"c", x"9", x"5", x"1", x"3", x"9", x"d", x"e", x"e", x"d", x"9", x"3", x"3", x"9", x"d", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"8", x"d", x"e", x"c", x"7", x"2", x"4", x"a", x"d", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"b", x"9", x"7", x"6", x"5", x"4", x"1", x"0", x"1", x"2", x"3", x"6", x"a", x"d", x"e", x"e", x"e", x"d", x"9", x"3", x"3", x"9", x"d", x"e", x"f", x"e", x"c", x"7", x"2", x"1", x"7", x"d", x"e", x"e", x"c", x"7", x"1", x"4", x"a", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"9", x"5", x"8", x"c", x"d", x"b", x"7", x"2", x"2", x"8", x"c", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"c", x"7", x"3", x"1", x"0", x"2", x"5", x"6", x"7", x"6", x"3", x"1", x"2", x"6", x"b", x"e", x"e", x"e", x"e", x"a", x"4", x"2", x"9", x"d", x"e", x"f", x"e", x"e", x"9", x"4", x"1", x"5", x"c", x"e", x"e", x"c", x"6", x"1", x"5", x"b", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"8", x"3", x"6", x"9", x"8", x"7", x"4", x"1", x"1", x"5", x"b", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"c", x"7", x"4", x"1", x"1", x"5", x"a", x"c", x"c", x"b", x"8", x"4", x"1", x"3", x"9", x"d", x"e", x"e", x"e", x"a", x"4", x"1", x"8", x"d", x"e", x"f", x"f", x"e", x"b", x"5", x"1", x"5", x"b", x"e", x"e", x"b", x"5", x"1", x"6", x"c", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"c", x"6", x"1", x"2", x"3", x"2", x"1", x"2", x"2", x"0", x"3", x"a", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"b", x"9", x"4", x"2", x"7", x"c", x"e", x"e", x"e", x"c", x"7", x"2", x"2", x"6", x"c", x"e", x"f", x"e", x"a", x"4", x"2", x"8", x"d", x"e", x"f", x"f", x"e", x"b", x"5", x"2", x"5", x"b", x"e", x"e", x"b", x"4", x"2", x"6", x"c", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"a", x"4", x"1", x"3", x"5", x"7", x"8", x"8", x"6", x"2", x"1", x"8", x"d", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"b", x"5", x"2", x"7", x"c", x"e", x"f", x"f", x"e", x"a", x"4", x"1", x"5", x"b", x"e", x"f", x"e", x"a", x"3", x"3", x"8", x"d", x"e", x"f", x"f", x"e", x"c", x"6", x"2", x"5", x"b", x"e", x"e", x"b", x"5", x"2", x"6", x"c", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"9", x"4", x"7", x"a", x"b", x"c", x"d", x"d", x"a", x"5", x"1", x"6", x"b", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"2", x"7", x"c", x"e", x"f", x"f", x"e", x"c", x"5", x"1", x"4", x"a", x"e", x"e", x"e", x"a", x"3", x"2", x"8", x"d", x"e", x"f", x"f", x"e", x"b", x"6", x"2", x"5", x"c", x"e", x"e", x"b", x"5", x"1", x"6", x"b", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"7", x"5", x"a", x"d", x"e", x"e", x"e", x"e", x"b", x"6", x"1", x"3", x"8", x"c", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"5", x"1", x"7", x"c", x"e", x"f", x"f", x"e", x"c", x"6", x"2", x"4", x"a", x"e", x"e", x"e", x"a", x"4", x"2", x"8", x"d", x"e", x"f", x"f", x"e", x"b", x"5", x"2", x"6", x"c", x"e", x"e", x"b", x"6", x"1", x"5", x"b", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"e", x"f", x"e", x"b", x"5", x"6", x"b", x"e", x"e", x"f", x"e", x"c", x"9", x"4", x"0", x"0", x"4", x"a", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"5", x"1", x"7", x"c", x"e", x"f", x"f", x"e", x"c", x"7", x"2", x"5", x"a", x"e", x"e", x"e", x"a", x"5", x"2", x"8", x"d", x"f", x"f", x"f", x"e", x"b", x"4", x"2", x"7", x"c", x"e", x"e", x"c", x"7", x"2", x"4", x"9", x"d", x"e", x"f", x"f", x"f", x"e", x"e", x"e", x"d", x"e", x"e", x"d", x"a", x"4", x"5", x"9", x"c", x"e", x"e", x"d", x"a", x"5", x"1", x"1", x"3", x"5", x"a", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"5", x"2", x"7", x"c", x"e", x"f", x"f", x"e", x"c", x"7", x"2", x"5", x"a", x"e", x"f", x"e", x"a", x"4", x"2", x"8", x"d", x"f", x"f", x"e", x"d", x"9", x"4", x"3", x"8", x"d", x"e", x"e", x"d", x"9", x"3", x"2", x"7", x"b", x"e", x"e", x"e", x"e", x"e", x"c", x"a", x"a", x"d", x"e", x"b", x"6", x"2", x"2", x"6", x"b", x"e", x"e", x"d", x"a", x"6", x"7", x"8", x"9", x"b", x"d", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"1", x"7", x"c", x"e", x"f", x"f", x"e", x"c", x"7", x"2", x"4", x"a", x"e", x"f", x"e", x"a", x"4", x"2", x"8", x"d", x"e", x"f", x"e", x"d", x"8", x"2", x"5", x"a", x"e", x"f", x"e", x"e", x"b", x"6", x"0", x"4", x"8", x"b", x"c", x"d", x"c", x"a", x"8", x"5", x"8", x"d", x"d", x"9", x"3", x"1", x"2", x"5", x"b", x"e", x"f", x"e", x"c", x"b", x"c", x"d", x"e", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"0", x"7", x"c", x"e", x"f", x"f", x"e", x"c", x"6", x"2", x"6", x"b", x"e", x"f", x"e", x"b", x"4", x"2", x"8", x"d", x"e", x"f", x"e", x"b", x"5", x"2", x"7", x"c", x"e", x"f", x"f", x"e", x"d", x"9", x"3", x"1", x"3", x"6", x"8", x"8", x"7", x"5", x"4", x"5", x"9", x"d", x"d", x"9", x"6", x"7", x"9", x"b", x"d", x"e", x"f", x"e", x"e", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"0", x"7", x"c", x"e", x"f", x"f", x"e", x"b", x"6", x"2", x"7", x"c", x"e", x"e", x"e", x"b", x"5", x"2", x"8", x"d", x"e", x"e", x"b", x"7", x"3", x"5", x"a", x"d", x"e", x"f", x"f", x"e", x"e", x"c", x"8", x"4", x"2", x"2", x"2", x"3", x"3", x"5", x"7", x"a", x"c", x"e", x"e", x"d", x"c", x"d", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"0", x"7", x"c", x"e", x"f", x"f", x"e", x"a", x"4", x"3", x"8", x"d", x"e", x"f", x"e", x"a", x"5", x"1", x"7", x"c", x"d", x"b", x"7", x"3", x"3", x"8", x"c", x"e", x"f", x"f", x"f", x"f", x"e", x"e", x"c", x"a", x"8", x"7", x"6", x"7", x"8", x"a", x"c", x"d", x"e", x"e", x"e", x"e", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"0", x"7", x"c", x"e", x"f", x"e", x"c", x"8", x"2", x"4", x"a", x"e", x"e", x"e", x"d", x"a", x"4", x"0", x"5", x"8", x"8", x"6", x"3", x"4", x"8", x"c", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"d", x"d", x"c", x"c", x"c", x"d", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"0", x"7", x"c", x"e", x"e", x"d", x"a", x"5", x"2", x"7", x"c", x"e", x"e", x"d", x"a", x"6", x"2", x"0", x"1", x"2", x"2", x"3", x"5", x"8", x"c", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"e", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"1", x"7", x"c", x"e", x"d", x"b", x"6", x"3", x"5", x"a", x"d", x"e", x"e", x"c", x"7", x"2", x"2", x"3", x"4", x"5", x"7", x"9", x"b", x"d", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"b", x"6", x"1", x"5", x"a", x"b", x"9", x"6", x"3", x"6", x"9", x"d", x"e", x"f", x"e", x"c", x"7", x"6", x"7", x"9", x"a", x"b", x"c", x"d", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"a", x"5", x"0", x"2", x"5", x"5", x"3", x"3", x"5", x"9", x"c", x"e", x"f", x"f", x"e", x"d", x"c", x"c", x"d", x"d", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"9", x"5", x"2", x"0", x"0", x"2", x"3", x"5", x"7", x"a", x"d", x"e", x"e", x"f", x"f", x"f", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"c", x"7", x"3", x"4", x"5", x"7", x"8", x"9", x"b", x"c", x"d", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"d", x"a", x"9", x"a", x"b", x"c", x"d", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"e", x"e", x"e", x"e", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"0", x"0", x"0", x"1", x"1", x"1", x"2", x"2", x"2", x"3", x"3", x"3", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"0", x"0", x"0", x"1", x"1", x"1", x"2", x"2", x"2", x"3", x"3", x"3", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"f", x"f", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"0", x"0", x"0", x"1", x"1", x"1", x"2", x"2", x"2", x"3", x"3", x"3", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"f", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"4", x"4", x"4", x"5", x"5", x"5", x"6", x"6", x"6", x"7", x"7", x"7", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"f", x"0", x"0", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"4", x"4", x"4", x"5", x"5", x"5", x"6", x"6", x"6", x"7", x"7", x"7", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"f", x"f", x"f", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"4", x"4", x"4", x"5", x"5", x"5", x"6", x"6", x"6", x"7", x"7", x"7", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"8", x"8", x"8", x"9", x"9", x"9", x"a", x"a", x"a", x"b", x"b", x"b", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"8", x"8", x"8", x"9", x"9", x"9", x"a", x"a", x"a", x"b", x"b", x"b", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"0", x"0", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"8", x"8", x"8", x"9", x"9", x"9", x"a", x"a", x"a", x"b", x"b", x"b", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"f", x"f", x"f", x"f", x"0", x"f", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"c", x"c", x"d", x"d", x"d", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"c", x"c", x"d", x"d", x"d", x"e", x"e", x"e", x"f", x"f", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"0", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"c", x"c", x"c", x"d", x"d", x"d", x"e", x"e", x"e", x"f", x"f", x"f", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"0", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f",
	x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f", x"f"
);
end package;
